module generate_round_keys(input wire clk, n_rst, input wire [63:0] key, input wire[1:0] mode, 
			   output wire[47:0] round1,round2,round3,round4,round5,round6,round7,round8,round9,round10,round11,round12,round13,round14,round15, round16);
	wire[27:0] l1,l2,l3,l4,l5,l6,l7,l8,l9,l10,l11,l12,l13,l14,l15,l16,
		r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16;
	wire[55:0] p, p1, p2, p3, p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,p16;
	wire [47:0] pp1,pp2,pp3,pp4,pp5,pp6,pp7,pp8,pp9,pp10,pp11,pp12,pp13,pp14,pp15,pp16;
	assign p[55:48] = {key[56],key[48],key[40],key[32],key[24],key[16],key[8],key[0]};
	assign p[47:40] = {key[57],key[49],key[41],key[33],key[25],key[17],key[9],key[1]};
	assign p[39:32] = {key[58],key[50],key[42],key[34],key[26],key[18],key[10],key[2]};
	assign p[31:24] = {key[59],key[51],key[43],key[35],key[62],key[54],key[46],key[38]};
	assign p[23:16] = {key[30],key[22],key[14],key[6],key[61],key[53],key[45],key[37]};
	assign p[15:8]  = {key[29],key[21],key[13],key[5],key[60],key[52],key[44],key[36]};
	assign p[7:0]   = {key[28],key[20],key[12],key[4],key[27],key[19],key[11],key[3]};
	assign l1	 = {p[26:0],p[27]};		//left shift 1
	assign r1 	 = {p[54:28],p[55]};		//left shift 1
	assign l2	 = {l1[26:0],l1[27]};	
	assign r2	 = {r1[26:0],r1[27]};
	assign l3	 = {l2[25:0], l2[27:26]};
	assign r3	 = {r2[25:0], r2[27:26]};
	assign l4	 = {l3[25:0], l3[27:26]};
	assign r4	 = {r3[25:0], r3[27:26]};
	assign l5	 = {l4[25:0], l4[27:26]};
	assign r5	 = {r4[25:0], r4[27:26]};
	assign l6	 = {l5[25:0], l5[27:26]};
	assign r6	 = {r5[25:0], r5[27:26]};
	assign l7	 = {l6[25:0], l6[27:26]};
	assign r7	 = {r6[25:0], r6[27:26]};
	assign l8	 = {l7[25:0], l7[27:26]};
	assign r8	 = {r7[25:0], r7[27:26]};
	assign l9	 = {l8[26:0],l8[27]};
	assign r9 	 = {r8[26:0],r8[27]};
	assign l10	 = {l9[25:0], l9[27:26]};
	assign r10	 = {r9[25:0], r9[27:26]};
	assign l11	 = {l10[25:0], l10[27:26]};
	assign r11	 = {r10[25:0], r10[27:26]};
	assign l12	 = {l11[25:0], l11[27:26]};
	assign r12	 = {r11[25:0], r11[27:26]};
	assign l13	 = {l12[25:0], l12[27:26]};
	assign r13	 = {r12[25:0], r12[27:26]};
	assign l14	 = {l13[25:0], l13[27:26]};
	assign r14	 = {r13[25:0], r13[27:26]};
	assign l15	 = {l14[25:0], l14[27:26]};
	assign r15	 = {r14[25:0], r14[27:26]};
	assign l16	 = {l15[26:0],l15[27]};
	assign r16 	 = {r15[26:0],r15[27]};
	assign p1	 = {r1, l1};
	assign p2	 = {r2, l2};
	assign p3	 = {r3, l3};
	assign p4	 = {r4, l4};
	assign p5	 = {r5, l5};
	assign p6	 = {r6, l6};
	assign p7	 = {r7, l7};
	assign p8	 = {r8, l8};
	assign p9	 = {r9, l9};
	assign p10	 = {r10, l10};
	assign p11	 = {r11, l11};
	assign p12	 = {r12, l12};
	assign p13	 = {r13, l13};
	assign p14	 = {r14, l14};
	assign p15	 = {r15, l15};
	assign p16	 = {r16, l16};
	assign pp1[47:40]	 = {p1[13],p1[16],p1[10],p1[23],p1[0],p1[4],p1[2],p1[27]};
	assign pp1[39:32]	 = {p1[14],p1[5],p1[20],p1[9],p1[22],p1[18],p1[11],p1[3]};
	assign pp1[31:24]	 = {p1[25],p1[7],p1[15],p1[6],p1[26],p1[19],p1[12],p1[1]};
	assign pp1[23:16]	 = {p1[40],p1[51],p1[30],p1[36],p1[46],p1[54],p1[29],p1[39]};
	assign pp1[15:8]	 = {p1[50],p1[44],p1[32],p1[47],p1[43],p1[48],p1[38],p1[55]};
	assign pp1[7:0]	 	 = {p1[33],p1[52],p1[45],p1[41],p1[49],p1[35],p1[28],p1[31]};

	assign pp2[47:40]	 = {p2[13],p2[16],p2[10],p2[23],p2[0],p2[4],p2[2],p2[27]};
	assign pp2[39:32]	 = {p2[14],p2[5],p2[20],p2[9],p2[22],p2[18],p2[11],p2[3]};
	assign pp2[31:24]	 = {p2[25],p2[7],p2[15],p2[6],p2[26],p2[19],p2[12],p2[1]};
	assign pp2[23:16]	 = {p2[40],p2[51],p2[30],p2[36],p2[46],p2[54],p2[29],p2[39]};
	assign pp2[15:8]	 = {p2[50],p2[44],p2[32],p2[47],p2[43],p2[48],p2[38],p2[55]};
	assign pp2[7:0]	 	 = {p2[33],p2[52],p2[45],p2[41],p2[49],p2[35],p2[28],p2[31]};

	assign pp3[47:40]	 = {p3[13],p3[16],p3[10],p3[23],p3[0],p3[4],p3[2],p3[27]};
	assign pp3[39:32]	 = {p3[14],p3[5],p3[20],p3[9],p3[22],p3[18],p3[11],p3[3]};
	assign pp3[31:24]	 = {p3[25],p3[7],p3[15],p3[6],p3[26],p3[19],p3[12],p3[1]};
	assign pp3[23:16]	 = {p3[40],p3[51],p3[30],p3[36],p3[46],p3[54],p3[29],p3[39]};
	assign pp3[15:8]	 = {p3[50],p3[44],p3[32],p3[47],p3[43],p3[48],p3[38],p3[55]};
	assign pp3[7:0]	 	 = {p3[33],p3[52],p3[45],p3[41],p3[49],p3[35],p3[28],p3[31]};

	assign pp4[47:40]	 = {p4[13],p4[16],p4[10],p4[23],p4[0],p4[4],p4[2],p4[27]};
	assign pp4[39:32]	 = {p4[14],p4[5],p4[20],p4[9],p4[22],p4[18],p4[11],p4[3]};
	assign pp4[31:24]	 = {p4[25],p4[7],p4[15],p4[6],p4[26],p4[19],p4[12],p4[1]};
	assign pp4[23:16]	 = {p4[40],p4[51],p4[30],p4[36],p4[46],p4[54],p4[29],p4[39]};
	assign pp4[15:8]	 = {p4[50],p4[44],p4[32],p4[47],p4[43],p4[48],p4[38],p4[55]};
	assign pp4[7:0]	 	 = {p4[33],p4[52],p4[45],p4[41],p4[49],p4[35],p4[28],p4[31]};

	assign pp5[47:40]	 = {p5[13],p5[16],p5[10],p5[23],p5[0],p5[4],p5[2],p5[27]};
	assign pp5[39:32]	 = {p5[14],p5[5],p5[20],p5[9],p5[22],p5[18],p5[11],p5[3]};
	assign pp5[31:24]	 = {p5[25],p5[7],p5[15],p5[6],p5[26],p5[19],p5[12],p5[1]};
	assign pp5[23:16]	 = {p5[40],p5[51],p5[30],p5[36],p5[46],p5[54],p5[29],p5[39]};
	assign pp5[15:8]	 = {p5[50],p5[44],p5[32],p5[47],p5[43],p5[48],p5[38],p5[55]};
	assign pp5[7:0]	 	 = {p5[33],p5[52],p5[45],p5[41],p5[49],p5[35],p5[28],p5[31]};

	assign pp6[47:40]	 = {p6[13],p6[16],p6[10],p6[23],p6[0],p6[4],p6[2],p6[27]};
	assign pp6[39:32]	 = {p6[14],p6[5],p6[20],p6[9],p6[22],p6[18],p6[11],p6[3]};
	assign pp6[31:24]	 = {p6[25],p6[7],p6[15],p6[6],p6[26],p6[19],p6[12],p6[1]};
	assign pp6[23:16]	 = {p6[40],p6[51],p6[30],p6[36],p6[46],p6[54],p6[29],p6[39]};
	assign pp6[15:8]	 = {p6[50],p6[44],p6[32],p6[47],p6[43],p6[48],p6[38],p6[55]};
	assign pp6[7:0]	 	 = {p6[33],p6[52],p6[45],p6[41],p6[49],p6[35],p6[28],p6[31]};

	assign pp7[47:40]	 = {p7[13],p7[16],p7[10],p7[23],p7[0],p7[4],p7[2],p7[27]};
	assign pp7[39:32]	 = {p7[14],p7[5],p7[20],p7[9],p7[22],p7[18],p7[11],p7[3]};
	assign pp7[31:24]	 = {p7[25],p7[7],p7[15],p7[6],p7[26],p7[19],p7[12],p7[1]};
	assign pp7[23:16]	 = {p7[40],p7[51],p7[30],p7[36],p7[46],p7[54],p7[29],p7[39]};
	assign pp7[15:8]	 = {p7[50],p7[44],p7[32],p7[47],p7[43],p7[48],p7[38],p7[55]};
	assign pp7[7:0]	 	 = {p7[33],p7[52],p7[45],p7[41],p7[49],p7[35],p7[28],p7[31]};

	assign pp8[47:40]	 = {p8[13],p8[16],p8[10],p8[23],p8[0],p8[4],p8[2],p8[27]};
	assign pp8[39:32]	 = {p8[14],p8[5],p8[20],p8[9],p8[22],p8[18],p8[11],p8[3]};
	assign pp8[31:24]	 = {p8[25],p8[7],p8[15],p8[6],p8[26],p8[19],p8[12],p8[1]};
	assign pp8[23:16]	 = {p8[40],p8[51],p8[30],p8[36],p8[46],p8[54],p8[29],p8[39]};
	assign pp8[15:8]	 = {p8[50],p8[44],p8[32],p8[47],p8[43],p8[48],p8[38],p8[55]};
	assign pp8[7:0]	 	 = {p8[33],p8[52],p8[45],p8[41],p8[49],p8[35],p8[28],p8[31]};

	assign pp9[47:40]	 = {p9[13],p9[16],p9[10],p9[23],p9[0],p9[4],p9[2],p9[27]};
	assign pp9[39:32]	 = {p9[14],p9[5],p9[20],p9[9],p9[22],p9[18],p9[11],p9[3]};
	assign pp9[31:24]	 = {p9[25],p9[7],p9[15],p9[6],p9[26],p9[19],p9[12],p9[1]};
	assign pp9[23:16]	 = {p9[40],p9[51],p9[30],p9[36],p9[46],p9[54],p9[29],p9[39]};
	assign pp9[15:8]	 = {p9[50],p9[44],p9[32],p9[47],p9[43],p9[48],p9[38],p9[55]};
	assign pp9[7:0]	 	 = {p9[33],p9[52],p9[45],p9[41],p9[49],p9[35],p9[28],p9[31]};

	assign pp10[47:40]	 = {p10[13],p10[16],p10[10],p10[23],p10[0],p10[4],p10[2],p10[27]};
	assign pp10[39:32]	 = {p10[14],p10[5],p10[20],p10[9],p10[22],p10[18],p10[11],p10[3]};
	assign pp10[31:24]	 = {p10[25],p10[7],p10[15],p10[6],p10[26],p10[19],p10[12],p10[1]};
	assign pp10[23:16]	 = {p10[40],p10[51],p10[30],p10[36],p10[46],p10[54],p10[29],p10[39]};
	assign pp10[15:8]	 = {p10[50],p10[44],p10[32],p10[47],p10[43],p10[48],p10[38],p10[55]};
	assign pp10[7:0]	 = {p10[33],p10[52],p10[45],p10[41],p10[49],p10[35],p10[28],p10[31]};

	assign pp11[47:40]	 = {p11[13],p11[16],p11[10],p11[23],p11[0],p11[4],p11[2],p11[27]};
	assign pp11[39:32]	 = {p11[14],p11[5],p11[20],p11[9],p11[22],p11[18],p11[11],p11[3]};
	assign pp11[31:24]	 = {p11[25],p11[7],p11[15],p11[6],p11[26],p11[19],p11[12],p11[1]};
	assign pp11[23:16]	 = {p11[40],p11[51],p11[30],p11[36],p11[46],p11[54],p11[29],p11[39]};
	assign pp11[15:8]	 = {p11[50],p11[44],p11[32],p11[47],p11[43],p11[48],p11[38],p11[55]};
	assign pp11[7:0]	 = {p11[33],p11[52],p11[45],p11[41],p11[49],p11[35],p11[28],p11[31]};

	assign pp12[47:40]	 = {p12[13],p12[16],p12[10],p12[23],p12[0],p12[4],p12[2],p12[27]};
	assign pp12[39:32]	 = {p12[14],p12[5],p12[20],p12[9],p12[22],p12[18],p12[11],p12[3]};
	assign pp12[31:24]	 = {p12[25],p12[7],p12[15],p12[6],p12[26],p12[19],p12[12],p12[1]};
	assign pp12[23:16]	 = {p12[40],p12[51],p12[30],p12[36],p12[46],p12[54],p12[29],p12[39]};
	assign pp12[15:8]	 = {p12[50],p12[44],p12[32],p12[47],p12[43],p12[48],p12[38],p12[55]};
	assign pp12[7:0]	 = {p12[33],p12[52],p12[45],p12[41],p12[49],p12[35],p12[28],p12[31]};

	assign pp13[47:40]	 = {p13[13],p13[16],p13[10],p13[23],p13[0],p13[4],p13[2],p13[27]};
	assign pp13[39:32]	 = {p13[14],p13[5],p13[20],p13[9],p13[22],p13[18],p13[11],p13[3]};
	assign pp13[31:24]	 = {p13[25],p13[7],p13[15],p13[6],p13[26],p13[19],p13[12],p13[1]};
	assign pp13[23:16]	 = {p13[40],p13[51],p13[30],p13[36],p13[46],p13[54],p13[29],p13[39]};
	assign pp13[15:8]	 = {p13[50],p13[44],p13[32],p13[47],p13[43],p13[48],p13[38],p13[55]};
	assign pp13[7:0]	 = {p13[33],p13[52],p13[45],p13[41],p13[49],p13[35],p13[28],p13[31]};

	assign pp14[47:40]	 = {p14[13],p14[16],p14[10],p14[23],p14[0],p14[4],p14[2],p14[27]};
	assign pp14[39:32]	 = {p14[14],p14[5],p14[20],p14[9],p14[22],p14[18],p14[11],p14[3]};
	assign pp14[31:24]	 = {p14[25],p14[7],p14[15],p14[6],p14[26],p14[19],p14[12],p14[1]};
	assign pp14[23:16]	 = {p14[40],p14[51],p14[30],p14[36],p14[46],p14[54],p14[29],p14[39]};
	assign pp14[15:8]	 = {p14[50],p14[44],p14[32],p14[47],p14[43],p14[48],p14[38],p14[55]};
	assign pp14[7:0]	 = {p14[33],p14[52],p14[45],p14[41],p14[49],p14[35],p14[28],p14[31]};

	assign pp15[47:40]	 = {p15[13],p15[16],p15[10],p15[23],p15[0],p15[4],p15[2],p15[27]};
	assign pp15[39:32]	 = {p15[14],p15[5],p15[20],p15[9],p15[22],p15[18],p15[11],p15[3]};
	assign pp15[31:24]	 = {p15[25],p15[7],p15[15],p15[6],p15[26],p15[19],p15[12],p15[1]};
	assign pp15[23:16]	 = {p15[40],p15[51],p15[30],p15[36],p15[46],p15[54],p15[29],p15[39]};
	assign pp15[15:8]	 = {p15[50],p15[44],p15[32],p15[47],p15[43],p15[48],p15[38],p15[55]};
	assign pp15[7:0]	 = {p15[33],p15[52],p15[45],p15[41],p15[49],p15[35],p15[28],p15[31]};

	assign pp16[47:40]	 = {p16[13],p16[16],p16[10],p16[23],p16[0],p16[4],p16[2],p16[27]};
	assign pp16[39:32]	 = {p16[14],p16[5],p16[20],p16[9],p16[22],p16[18],p16[11],p16[3]};
	assign pp16[31:24]	 = {p16[25],p16[7],p16[15],p16[6],p16[26],p16[19],p16[12],p16[1]};
	assign pp16[23:16]	 = {p16[40],p16[51],p16[30],p16[36],p16[46],p16[54],p16[29],p16[39]};
	assign pp16[15:8]	 = {p16[50],p16[44],p16[32],p16[47],p16[43],p16[48],p16[38],p16[55]};
	assign pp16[7:0]	 = {p16[33],p16[52],p16[45],p16[41],p16[49],p16[35],p16[28],p16[31]};
	


	assign round1 = (mode == 2'b00) ? pp1 : (mode == 2'b01) ? pp16 : 48'd0;
	assign round2 = (mode == 2'b00) ? pp2 : (mode == 2'b01) ? pp15 : 48'd0;
	assign round3 = (mode == 2'b00) ? pp3 : (mode == 2'b01) ? pp14 : 48'd0;
	assign round4 = (mode == 2'b00) ? pp4 : (mode == 2'b01) ? pp13 : 48'd0;
	assign round5 = (mode == 2'b00) ? pp5 : (mode == 2'b01) ? pp12 : 48'd0;
	assign round6 = (mode == 2'b00) ? pp6 : (mode == 2'b01) ? pp11 : 48'd0;
	assign round7 = (mode == 2'b00) ? pp7 : (mode == 2'b01) ? pp10 : 48'd0;
	assign round8 = (mode == 2'b00) ? pp8 : (mode == 2'b01) ? pp9 : 48'd0;
	assign round9 = (mode == 2'b00) ? pp9 : (mode == 2'b01) ? pp8 : 48'd0;
	assign round10 = (mode == 2'b00) ? pp10 : (mode == 2'b01) ? pp7 : 48'd0;
	assign round11 = (mode == 2'b00) ? pp11 : (mode == 2'b01) ? pp6 : 48'd0;
	assign round12 = (mode == 2'b00) ? pp12 : (mode == 2'b01) ? pp5 : 48'd0;
	assign round13 = (mode == 2'b00) ? pp13 : (mode == 2'b01) ? pp4 : 48'd0;
	assign round14 = (mode == 2'b00) ? pp14 : (mode == 2'b01) ? pp3 : 48'd0;
	assign round15 = (mode == 2'b00) ? pp15 : (mode == 2'b01) ? pp2 : 48'd0;
	assign round16 = (mode == 2'b00) ? pp16 : (mode == 2'b01) ? pp1 : 48'd0;

endmodule
